// top

module top ( clk,
             rst,
			 // Instruction Memory
			 IM_Address,
             		 Instruction,
			 // Data Memory
			 DM_Address,
			 DM_enable,
			 DM_Write_Data,
			 DM_Read_Data);

	parameter data_size = 32;
	parameter mem_size = 16;
	parameter pc_size = 18;

	input  clk, rst;
	
	// Instruction Memory
	output [mem_size-1:0] IM_Address;	
	input  [data_size-1:0] Instruction;

	// Data Memory
	output [mem_size-1:0] DM_Address;
	output DM_enable;
	output [data_size-1:0] DM_Write_Data;	
    	input  [data_size-1:0] DM_Read_Data;
	
	// ALU
	wire [data_size-1:0] src2;
	wire [4:0] shamt;	
	wire [data_size-1:0] ALU_result;
	wire Zero;

	// Controller
	wire [5:0] opcode;
	wire [5:0] funct;
	wire [3:0] ALUOp;
	wire Reg_imm;
	wire RegWrite;
	wire MemtoReg;
	wire MemWrite;
	wire Branch;
	wire J;
	wire Jal;
	wire Jr;
	wire Half;

	// PC
	wire [pc_size-1:0] PCout;
	wire [pc_size-1:0] PC_add4;
	wire [pc_size-1:0] PC_add8;

	//Jump Part
	wire [pc_size-1:0] BranchAddr;
	wire [pc_size-1:0] JumpAddr;
	wire [1:0] JumpOP;
	wire [pc_size-1:0] PCin;
	
	// Regfile
	wire [4:0] Rd;
	wire [4:0] Rs;
	wire [4:0] Rt;
	wire [4:0] Rd_Rt_out;
	wire [4:0] WR_out;
	wire [data_size-1:0] WD_data;
	wire [data_size-1:0] WD_out;
	wire [data_size-1:0] Rs_data;
	wire [data_size-1:0] Rt_data;
	
	// Sign_extend	
	wire [15:0] imm;
	wire [data_size-1:0] imm_extend;

	// write back
	wire [data_size-1:0] WB_data;

	/* Wire connect-----------------------------------------------*/
	
	// ALU
	assign shamt = Instruction[10:6];
	assign JumpAddr = {Instruction[15:0],2'b0};

	// Controller
	assign opcode = Instruction[31:26];
	assign funct = Instruction[5:0];

	// PC
	assign IM_Address = PCout[pc_size-1:2];		

	// Registers
	assign Rd = Instruction[15:11];
	assign Rs = Instruction[25:21];
	assign Rt = Instruction[20:16];

	// Sign_extend
	assign imm = Instruction[15:0];
		
	// Data Memory
	assign DM_Address = ALU_result[17:2];
	assign DM_enable = MemWrite;
	assign DM_Write_Data = Rt_data;
	
	/* CPU---------------------------------------------------------*/
	
	// PC
	PC PC_component ( .clk(clk), .rst(rst), .PCin(PCin), .PCout(PCout));
					   
	ADD#(pc_size) ADD_Plus4 ( .A(PCout), .B(18'd4), .Cout(PC_add4));
	
	ADD#(pc_size) ADD_Plus_other_4 ( .A(PC_add4), .B(18'd4), .Cout(PC_add8));
	
	// Controller
	Controller Controller_component ( .opcode(opcode), .funct(funct), .ALUOp(ALUOp), .Reg_imm(Reg_imm), .RegWrite(RegWrite),
		.MemtoReg(MemtoReg), .MemWrite(MemWrite), .J(J), .Branch(Branch), .Jal(Jal), .Jr(Jr), .Half(Half));
	
	// Registers
	Mux2to1#(5) Rd_Rt ( .I0(Rd), .I1(Rt), .S(Reg_imm), .out(Rd_Rt_out));

	Mux2to1#(5) WR ( .I0(Rd_Rt_out), .I1(5'd31), .S(Jal), .out(WR_out));

	Mux2to1#(data_size) WD_Half ( .I0(WB_data),
		.I1({WB_data[15],WB_data[15],WB_data[15],WB_data[15],WB_data[15],WB_data[15],WB_data[15],WB_data[15],
			WB_data[15],WB_data[15],WB_data[15],WB_data[15],WB_data[15],WB_data[15],WB_data[15],WB_data[15],WB_data[15:0]}),
		.S(Half), .out(WD_data) );

	Mux2to1#(data_size) WD ( .I0(WD_data), .I1({14'b0,PC_add8}), .S(Jal), .out(WD_out));

	Regfile Regfile_component ( .clk(clk), .rst(rst), .Read_addr_1(Rs), .Read_addr_2(Rt), .Read_data_1(Rs_data), .Read_data_2(Rt_data),
		.RegWrite(RegWrite), .Write_addr(WR_out), .Write_data(WD_out));
	
	// sign_extend	
	Sign_extend extension ( .in(imm), .out(imm_extend));
	
	// ALU
	Mux2to1#(data_size) Rt_imm ( .I0(Rt_data), .I1(imm_extend), .S(Reg_imm), .out(src2));
	
	ALU ALU_component ( .ALUOp(ALUOp), .src1(Rs_data), .src2(src2), .shamt(shamt), .ALU_result(ALU_result), .Zero(Zero));
	
	//Jump Part
	ADD#(pc_size) ADD_Branch ( .A(PC_add4), .B({imm_extend[15:0],2'b0}), .Cout(BranchAddr));
	
	Jump_Ctrl Jump_Ctrl_component ( .Branch(Branch), .Zero(Zero), .Jr(Jr), .J(J), .JumpOP(JumpOP));

	Mux4to1 PC_Mux ( .I0(PC_add4), .I1(BranchAddr), .I2(Rs_data[pc_size-1:0]), .I3(JumpAddr), .S(JumpOP), .out(PCin));

	// write back
	Mux2to1#(data_size) WB_Mux ( .I0(ALU_result), .I1(DM_Read_Data), .S(MemtoReg), .out(WB_data));
	
endmodule





