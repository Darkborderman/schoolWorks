module rip_4bit(input1,input2,cin,sum,cout);

input [3:0]input1;
input [3:0]input2;
input cin;
output [3:0]sum;
output cout;


endmodule

