module F_adder(input1,input2,cin,sum,cout);

input input1,input2,cin;
output sum,cout;


endmodule

